// key scheduling